----------------------------------------------------------------------------------------
-- Archivo: bintobcd.vhd
----------------------------------------------------------------------------------------
-- Autor:     Mg. Ing. Mario Raffo
-- Email:     mraffo@pucp.edu.pe
-- Entidad:   Pontificia Universidad Católica del Perú (PUCP)
-- Facultad:  Estudios Generales Ciencias (EE.GG.CC) 
-- Curso:     1IEE04 - Diseño Digital
----------------------------------------------------------------------------------------
-- Historia de Versión:
-- Versión 1.0 (12/10/2017) - Mario Raffo 
----------------------------------------------------------------------------------------
-- Descripción:
-- Circuito que realiza un conversor de binario a bcd
----------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity bintobcd1 is
  port(signal a  :  in std_logic_vector(7 downto 0);
	   signal f  : out std_logic_vector(11 downto 0)) ;
end bintobcd1;

architecture structural of bintobcd1 is

  constant DONT_CARE : std_logic_vector(11 downto 0):= (others => '-');
  
  signal a_int : std_logic_vector(11 downto 0);

begin

  a_int <= "0000" & a;

  with a_int select
    f <= x"000" when x"000",
         x"001" when x"001",
         x"002" when x"002",
         x"003" when x"003",
         x"004" when x"004",
         x"005" when x"005",
         x"006" when x"006",
         x"007" when x"007",
         x"008" when x"008",
         x"009" when x"009",			 
         x"010" when x"00A",
         x"011" when x"00b",
         x"012" when x"00C",
         x"013" when x"00d",
         x"014" when x"00E",
         x"015" when x"00F",
         x"016" when x"010",
         x"017" when x"011",		 
         x"018" when x"012",
         x"019" when x"013",
         x"020" when x"014",	
         x"021" when x"015",
         x"022" when x"016",		 
         x"023" when x"017",
         x"024" when x"018",
         x"025" when x"019",	
         x"026" when x"01A",
         x"027" when x"01b",		 
         x"028" when x"01C",
         x"029" when x"01d",
         x"030" when x"01E",	
         x"031" when x"01F",	 
         x"032" when x"020",
         x"033" when x"021",
         x"034" when x"022",
         x"035" when x"023",
         x"036" when x"024",
         x"037" when x"025",
         x"038" when x"026",
         x"039" when x"027",
         x"040" when x"028",
         x"041" when x"029",			 
         x"042" when x"02A",
         x"043" when x"02b",
         x"044" when x"02C",
         x"045" when x"02d",
         x"046" when x"02E",
         x"047" when x"02F",
         x"048" when x"030",
         x"049" when x"031",		 
         x"050" when x"032",
         x"051" when x"033",
         x"052" when x"034",	
         x"053" when x"035",
         x"054" when x"036",		 
         x"055" when x"037",
         x"056" when x"038",
         x"057" when x"039",	
         x"058" when x"03A",
         x"059" when x"03b",		 
         x"060" when x"03C",
         x"061" when x"03D",
         x"062" when x"03E",	
         x"063" when x"03F",
			x"064" when x"040",
			x"065" when x"041",
         x"066" when x"042",
         x"067" when x"043",
         x"068" when x"044",
         x"069" when x"045",
         x"070" when x"046",
         x"071" when x"047",
         x"072" when x"048",
         x"073" when x"049",			 
         x"074" when x"04A",
         x"075" when x"04b",
         x"076" when x"04C",
         x"077" when x"04d",
         x"078" when x"04E",
         x"079" when x"04F",
         x"080" when x"050",
         x"081" when x"051",		 
         x"082" when x"052",
         x"083" when x"053",
         x"084" when x"054",	
         x"085" when x"055",
         x"086" when x"056",		 
         x"087" when x"057",
         x"088" when x"058",
         x"089" when x"059",	
         x"090" when x"05A",
         x"091" when x"05b",		 
         x"092" when x"05C",
         x"093" when x"05d",
         x"094" when x"05E",	
         x"095" when x"05F",	 
         x"096" when x"060",
         x"097" when x"061",
         x"098" when x"062",
         x"099" when x"063",
         x"100" when x"064",
         x"101" when x"065",
         x"102" when x"066",
         x"103" when x"067",
         x"104" when x"068",
         x"105" when x"069",			 
         x"106" when x"06A",
         x"107" when x"06b",
         x"108" when x"06C",
         x"109" when x"06d",
         x"110" when x"06E",
         x"111" when x"06F",
         x"112" when x"070",
         x"113" when x"071",		 
         x"114" when x"072",
         x"115" when x"073",
         x"116" when x"074",	
         x"117" when x"075",
         x"118" when x"076",		 
         x"119" when x"077",
         x"120" when x"078",
         x"121" when x"079",	
         x"122" when x"07A",
         x"123" when x"07b",		 
         x"124" when x"07C",
         x"125" when x"07D",
         x"126" when x"07E",	
         x"127" when x"07F",
			x"128" when x"080",
         x"129" when x"081",
         x"130" when x"082",	
         x"131" when x"083",	 
         x"132" when x"084",
         x"133" when x"085",
         x"134" when x"086",
         x"135" when x"087",
         x"136" when x"088",
         x"137" when x"089",
         x"138" when x"08A",
         x"139" when x"08B",
         x"140" when x"08C",
         x"141" when x"08D",			 
         x"142" when x"08E",
         x"143" when x"08F",
         x"144" when x"090",
         x"145" when x"091",
         x"146" when x"092",
         x"147" when x"093",
         x"148" when x"094",
         x"149" when x"095",		 
         x"150" when x"096",
         x"151" when x"097",
         x"152" when x"098",	
         x"153" when x"099",
         x"154" when x"09A",		 
         x"155" when x"09B",
         x"156" when x"09C",
         x"157" when x"09d",	
         x"158" when x"09e",
         x"159" when x"09f",		 
         x"160" when x"0a0",
         x"161" when x"0a1",
         x"162" when x"0a2",	
         x"163" when x"0a3",
			x"164" when x"0a4",
			x"165" when x"0a5",
         x"166" when x"0a6",
         x"167" when x"0a7",
         x"168" when x"0a8",
         x"169" when x"0a9",
         x"170" when x"0aa",
         x"171" when x"0ab",
         x"172" when x"0ac",
         x"173" when x"0ad",			 
         x"174" when x"0ae",
         x"175" when x"0af",
         x"176" when x"0b0",
         x"177" when x"0b1",
         x"178" when x"0b2",
         x"179" when x"0b3",
         x"180" when x"0b4",
         x"181" when x"0b5",		 
         x"182" when x"0b6",
         x"183" when x"0b7",
         x"184" when x"0b8",	
         x"185" when x"0b9",
         x"186" when x"0ba",		 
         x"187" when x"0bb",
         x"188" when x"0bc",
         x"189" when x"0bd",	
         x"190" when x"0be",
         x"191" when x"0bf",		 
         x"192" when x"0c0",
         x"193" when x"0c1",
         x"194" when x"0c2",	
         x"195" when x"0c3",	 
         x"196" when x"0c4",
         x"197" when x"0c5",
         x"198" when x"0c6",
         x"199" when x"0c7",
			x"200" when x"0c8",
         x"201" when x"0c9",
         x"202" when x"0ca",
         x"203" when x"0cb",
         x"204" when x"0cc",
         x"205" when x"0cd",
         x"206" when x"0ce",
         x"207" when x"0cf",
         x"208" when x"0d0",
         x"209" when x"0d1",			 
         x"210" when x"0d2",
         x"211" when x"0d3",
         x"212" when x"0d4",
         x"213" when x"0d5",
         x"214" when x"0d6",
         x"215" when x"0d7",
         x"216" when x"0d8",
         x"217" when x"0d9",		 
         x"218" when x"0da",
         x"219" when x"0db",
         x"220" when x"0dc",	
         x"221" when x"0dd",
         x"222" when x"0de",		 
         x"223" when x"0df",
         x"224" when x"0e0",
         x"225" when x"0e1",	
         x"226" when x"0e2",
         x"227" when x"0e3",		 
         x"228" when x"0e4",
         x"229" when x"0e5",
         x"230" when x"0e6",	
         x"231" when x"0e7",	 
         x"232" when x"0e8",
         x"233" when x"0e9",
         x"234" when x"0ea",
         x"235" when x"0eb",
         x"236" when x"0ec",
         x"237" when x"0ed",
         x"238" when x"0ee",
         x"239" when x"0ef",
         x"240" when x"0f0",
         x"241" when x"0f1",			 
         x"242" when x"0f2",
         x"243" when x"0f3",
         x"244" when x"0f4",
         x"245" when x"0f5",
         x"246" when x"0f6",
         x"247" when x"0f7",
         x"248" when x"0f8",
         x"249" when x"0f9",		 
         x"250" when x"0fa",
         x"251" when x"0fb",
         x"252" when x"0fc",	
         x"253" when x"0fd",
         x"254" when x"0fe",		 
         x"255" when x"0ff",
         DONT_CARE when others;

end structural;